`timescale 1ns / 1ps
module alu_tb();
    reg signed [31:0]a,b;
    reg [3:0]sel;
    wire signed [31:0]out;
    wire signed [63:0] out_m;
    wire zf,cf,nf,of;
    signed_controller c1(a,b,sel,out,out_m,cf,zf,of,nf);
    initial begin
        a=32'sd777965536;b=-32'sd687544332;sel=4'b0000;//and gate
        #10 a=32'sd430965904;b=32'sd4357764;
        #10 a=-32'sd5609545;b=-32'sd4690590;
        #10 a=32'sd777965536;b=-32'sd687544332;sel=4'b0001;//or gate
        #10 a=32'sd430965904;b=32'sd4357764;
        #10 a=-32'sd5609545;b=-32'sd4690590;
        #10 a=32'sd777965536;b=-32'sd687544332;sel=4'b0010;//xor gate
        #10 a=32'sd430965904;b=32'sd4357764;
        #10 a=-32'sd5609545;b=-32'sd4690590;
        #10 a=32'sd777965536;b=-32'sd687544332;sel=4'b0011;//not gate
        #10 a=32'sd430965904;b=32'sd4357764;
        #10 a=-32'sd5609545;b=-32'sd4690590;
        #10 a=32'sd777965536;b=-32'sd987544332;sel=4'b0100;//add
        #10 a=32'sd430965904;b=-32'sd4357764;
        #10 a=-32'sd5609545;b=-32'sd4690590;
        #10 a=32'sd564398597;b=32'sd968439569;
        #10 a=32'sd496569044;b=-32'sd496569044;
        #10 a=32'sd1973741829;b=32'sd1973741829;
        #10 a=32'sd777965536;b=-32'sd987544332;sel=4'b0101;//sub
        #10 a=32'sd430965904;b=-32'sd4357764;
        #10 a=-32'sd5609545;b=-32'sd4690590;
        #10 a=32'sd564398597;b=32'sd968439569;
        #10 a=32'sd496569044;b=32'sd496569044;
        #10 a=-32'sd1973741829;b=32'sd1973741829;
        #10 a=32'sd777965536;b=-32'sd987544332;sel=4'b0110;//mul
        #10 a=32'sd430965904;b=-32'sd4357764;
        #10 a=-32'sd5609545;b=-32'sd4690590;
        #10 a=32'sd564398597;b=32'sd968439569;
        #10 a=32'sd496569044;b=-32'sd496569044;
        #10 a=32'sd329373247;b=5'd12;sel=4'b0111;//arithmetic right shift
        #10 a=-32'sd893483234;b=5'd23;sel=4'b1000;//left shift
        #10 a=32'sd1973741829;b=5'd1;
        #10 a=32'sd43932754;b=5'd31;
        #10 a=-32'd32653565;b=5'd31;sel=4'b0111;
        #10 a=32'sd5398457;b=32'sd90505443;sel=4'b1001;//less than
        #10 a=-32'sd4096580;b=32'sd0956445;sel=4'b1010;//equal
        #10 a=32'sd436907954;b=-32'sd497843978;sel=4'b1011;//greter than
        #10 a=-32'sd43984379;b=-32'sd43984379;sel=4'b1010;//equal
        #10 a=-32'sd90319842;b=-32'sd28648976;sel=4'b1111;//default
        #10 $finish;
    end
    initial 
        $monitor("%g %sb %sb %b %sb %sb %b %b %b %b",$time,a,b,sel,out,out_m,zf,cf,nf,of);
endmodule